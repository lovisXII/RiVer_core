import riscv::*;

module rename (
)
endmodule