// This module must instanciate the interface between the fetch unit and the caches
// It can fetch several instruction at the same cycle so it must be parametrizable