import riscv::*;

module arith_queue(
    input logic instr,
    output logic issue_instr,
)
endmodule