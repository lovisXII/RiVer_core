module decoder import riscv_pkg::*;(
    input logic[XLEN-1:0] instr_i;
    input logic[XLEN-1:0] pc_i;
);



endmodule